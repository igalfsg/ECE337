// $Id: $
// File name:   moor.sv
// Created:     2/4/2016
// Author:      Igal Flegmann Sandler
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: first lab thing.
